// Copyright (c) 2014-2025 John Seamons, ZL4VO/KF6VO

`timescale 1ns / 100ps

module IQ_SAMPLER_4K_32B ();
        
endmodule
