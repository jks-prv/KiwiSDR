localparam RX_CFG = 44;
`define USE_WF
